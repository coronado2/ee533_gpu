// 8 registers x 64-bit. Uses two BRAM instances mirrored for 2R/1W.

module regfile_bram (
    input  wire        clk,

    // Read port A (rs1)
    input  wire [2:0]  rs1_addr,
    output wire [63:0] rs1_data,

    // Read port B (rs2)
    input  wire [2:0]  rs2_addr,
    output wire [63:0] rs2_data,

    // Write port
    input  wire        we,
    input  wire [2:0]  rd_addr,
    input  wire [63:0] rd_data
);

// --- BRAM A (for rs1 read) ---
// Connect to Block Memory Generator IP instance "regfile_bram0"
// Ports naming below are typical; adjust per IP wrapper generated by Vivado.
// This is a template connection: update port names to match your IP instance.

regfile_bram0 u_bram0 (
    .clka(clk),
    .ena(1'b1),
    .wea(we),
    .addra(rd_addr), // write address (write-first behavior recommended)
    .dina(rd_data),
    .douta(),        // unused

    .clkb(clk),
    .enb(1'b1),
    .web(1'b0),
    .addrb(rs1_addr),
    .dinb(64'd0),
    .doutb(rs1_data)
);

// --- BRAM B (for rs2 read) ---
// Connect to Block Memory Generator IP instance "regfile_bram1"
regfile_bram1 u_bram1 (
    .clka(clk),
    .ena(1'b1),
    .wea(we),
    .addra(rd_addr), // write address (mirror write)
    .dina(rd_data),
    .douta(), 

    .clkb(clk),
    .enb(1'b1),
    .web(1'b0),
    .addrb(rs2_addr),
    .dinb(64'd0),
    .doutb(rs2_data)
);

endmodule
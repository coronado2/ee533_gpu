// tensor_bf16_4lane.v  (full version)
//
// 4-lane BFloat16 tensor unit supporting:
//   OP_VADD  (3'b000) ? element-wise addition:       rd = a + b
//   OP_VSUB  (3'b001) ? element-wise subtraction:    rd = a - b
//   OP_VMUL  (3'b010) ? element-wise multiply:       rd = a * b
//   OP_FMAC  (3'b011) ? fused multiply-accumulate:   rd = a * b + acc
//   OP_RELU  (3'b100) ? ReLU on a:                   rd = max(0, a)
//
// Each 64-bit register holds 4 packed BF16 values:
//   lane0=[15:0], lane1=[31:16], lane2=[47:32], lane3=[63:48]
//
// Latency by operation:
//   VADD / VSUB : 3 cycles  (bf16_add latency)
//   VMUL        : 2 cycles  (bf16_mul latency)
//   FMAC        : 5 cycles  (mul=2, add=3 chained)
//   RELU        : 1 cycle   (combinational + 1 reg stage)
//
// Interface:
//   start  ? assert for 1 cycle to latch inputs and begin
//   op     ? operation select (held stable until done)
//   done   ? pulses high for exactly 1 cycle when rd_reg is valid

`define OP_VADD 3'b000
`define OP_VSUB 3'b001
`define OP_VMUL 3'b010
`define OP_FMAC 3'b011
`define OP_RELU 3'b100

module tensor (
    input  wire        clk,
    input  wire        rst_n,
    input  wire        start,
    input  wire [2:0]  op,       // operation select
    input  wire [63:0] a_reg,    // packed 4x bf16
    input  wire [63:0] b_reg,    // packed 4x bf16
    input  wire [63:0] acc_reg,  // packed 4x bf16 accumulator (used by FMAC)
    output reg  [63:0] rd_reg,   // packed 4x bf16 result
    output reg         done
);

// ?????????????????????????????????????????????????????????????????????????????
// Unpack lanes
// ?????????????????????????????????????????????????????????????????????????????
wire [15:0] a0 = a_reg[15:0];  wire [15:0] a1 = a_reg[31:16];
wire [15:0] a2 = a_reg[47:32]; wire [15:0] a3 = a_reg[63:48];

wire [15:0] b0 = b_reg[15:0];  wire [15:0] b1 = b_reg[31:16];
wire [15:0] b2 = b_reg[47:32]; wire [15:0] b3 = b_reg[63:48];

wire [15:0] acc0 = acc_reg[15:0];  wire [15:0] acc1 = acc_reg[31:16];
wire [15:0] acc2 = acc_reg[47:32]; wire [15:0] acc3 = acc_reg[63:48];

// ?????????????????????????????????????????????????????????????????????????????
// Latch inputs on start (prevents glitches during multi-cycle ops)
// ?????????????????????????????????????????????????????????????????????????????
reg [63:0] a_lat, b_lat, acc_lat;
reg [2:0]  op_lat;
reg        running;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        a_lat   <= 64'd0;
        b_lat   <= 64'd0;
        acc_lat <= 64'd0;
        op_lat  <= 3'd0;
        running <= 1'b0;
    end else begin
        if (start) begin
            a_lat   <= a_reg;
            b_lat   <= b_reg;
            acc_lat <= acc_reg;
            op_lat  <= op;
            running <= 1'b1;
        end
        if (done) running <= 1'b0;
    end
end

// ?????????????????????????????????????????????????????????????????????????????
// OP_VADD / OP_VSUB  ? direct adder launch
// For subtraction we flip the sign bit of b before feeding bf16_add
// ?????????????????????????????????????????????????????????????????????????????
wire start_add = start && ((op == `OP_VADD) || (op == `OP_VSUB));

// B operand sign-flipped for subtraction
wire [15:0] b0_eff = (op == `OP_VSUB) ? {~b0[15], b0[14:0]} : b0;
wire [15:0] b1_eff = (op == `OP_VSUB) ? {~b1[15], b1[14:0]} : b1;
wire [15:0] b2_eff = (op == `OP_VSUB) ? {~b2[15], b2[14:0]} : b2;
wire [15:0] b3_eff = (op == `OP_VSUB) ? {~b3[15], b3[14:0]} : b3;

wire [15:0] addAB0_out, addAB1_out, addAB2_out, addAB3_out;
wire        addAB0_done, addAB1_done, addAB2_done, addAB3_done;

bf16_add u_addAB0 (.clk(clk), .rst_n(rst_n), .start(start_add),
                   .a(a0), .b(b0_eff), .y(addAB0_out), .done(addAB0_done));
bf16_add u_addAB1 (.clk(clk), .rst_n(rst_n), .start(start_add),
                   .a(a1), .b(b1_eff), .y(addAB1_out), .done(addAB1_done));
bf16_add u_addAB2 (.clk(clk), .rst_n(rst_n), .start(start_add),
                   .a(a2), .b(b2_eff), .y(addAB2_out), .done(addAB2_done));
bf16_add u_addAB3 (.clk(clk), .rst_n(rst_n), .start(start_add),
                   .a(a3), .b(b3_eff), .y(addAB3_out), .done(addAB3_done));

// ?????????????????????????????????????????????????????????????????????????????
// OP_VMUL ? multipliers only
// ?????????????????????????????????????????????????????????????????????????????
wire start_mul_direct = start && (op == `OP_VMUL);
// FMAC also needs multipliers (shares the same instances ? gated by start signal)
wire start_mul_fmac   = start && (op == `OP_FMAC);
wire start_mul = start_mul_direct | start_mul_fmac;

wire [15:0] mul0_out, mul1_out, mul2_out, mul3_out;
wire        mul0_done, mul1_done, mul2_done, mul3_done;

bf16_mul u_mul0 (.clk(clk), .rst_n(rst_n), .start(start_mul),
                 .a(a0), .b(b0), .y(mul0_out), .done(mul0_done));
bf16_mul u_mul1 (.clk(clk), .rst_n(rst_n), .start(start_mul),
                 .a(a1), .b(b1), .y(mul1_out), .done(mul1_done));
bf16_mul u_mul2 (.clk(clk), .rst_n(rst_n), .start(start_mul),
                 .a(a2), .b(b2), .y(mul2_out), .done(mul2_done));
bf16_mul u_mul3 (.clk(clk), .rst_n(rst_n), .start(start_mul),
                 .a(a3), .b(b3), .y(mul3_out), .done(mul3_done));

// ?????????????????????????????????????????????????????????????????????????????
// OP_FMAC ? adder stage chained after multipliers (uses mul*_done as start)
// Only fire if op_lat is FMAC so the adders don't misfire on plain VMUL
// ?????????????????????????????????????????????????????????????????????????????
wire fmac_add_start0 = mul0_done && (op_lat == `OP_FMAC);
wire fmac_add_start1 = mul1_done && (op_lat == `OP_FMAC);
wire fmac_add_start2 = mul2_done && (op_lat == `OP_FMAC);
wire fmac_add_start3 = mul3_done && (op_lat == `OP_FMAC);

wire [15:0] add0_out, add1_out, add2_out, add3_out;
wire        add0_done, add1_done, add2_done, add3_done;

bf16_add u_add0 (.clk(clk), .rst_n(rst_n), .start(fmac_add_start0),
                 .a(acc_lat[15:0]),  .b(mul0_out), .y(add0_out), .done(add0_done));
bf16_add u_add1 (.clk(clk), .rst_n(rst_n), .start(fmac_add_start1),
                 .a(acc_lat[31:16]), .b(mul1_out), .y(add1_out), .done(add1_done));
bf16_add u_add2 (.clk(clk), .rst_n(rst_n), .start(fmac_add_start2),
                 .a(acc_lat[47:32]), .b(mul2_out), .y(add2_out), .done(add2_done));
bf16_add u_add3 (.clk(clk), .rst_n(rst_n), .start(fmac_add_start3),
                 .a(acc_lat[63:48]), .b(mul3_out), .y(add3_out), .done(add3_done));

// ?????????????????????????????????????????????????????????????????????????????
// OP_RELU ? combinational, registered 1 cycle after start
// ReLU: if sign bit is 1 (negative) ? output 0; else pass through.
// BF16 zero = 16'h0000.  Works for �0 correctly.
// ?????????????????????????????????????????????????????????????????????????????
wire [15:0] relu0 = a0[15] ? 16'h0000 : a0;
wire [15:0] relu1 = a1[15] ? 16'h0000 : a1;
wire [15:0] relu2 = a2[15] ? 16'h0000 : a2;
wire [15:0] relu3 = a3[15] ? 16'h0000 : a3;

reg [63:0] relu_result;
reg        relu_done;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        relu_result <= 64'd0;
        relu_done   <= 1'b0;
    end else begin
        relu_done <= (start && (op == `OP_RELU));
        if (start && (op == `OP_RELU))
            relu_result <= {relu3, relu2, relu1, relu0};
    end
end

// ?????????????????????????????????????????????????????????????????????????????
// Output mux ? select result based on latched op
// ?????????????????????????????????????????????????????????????????????????????
wire vadd_done = addAB0_done & addAB1_done & addAB2_done & addAB3_done
                 && (op_lat == `OP_VADD || op_lat == `OP_VSUB);

wire vmul_done = mul0_done & mul1_done & mul2_done & mul3_done
                 && (op_lat == `OP_VMUL);

wire fmac_done = add0_done & add1_done & add2_done & add3_done
                 && (op_lat == `OP_FMAC);

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        rd_reg <= 64'd0;
        done   <= 1'b0;
    end else begin
        done <= 1'b0; // default de-assert

        if (vadd_done) begin
            rd_reg <= {addAB3_out, addAB2_out, addAB1_out, addAB0_out};
            done   <= 1'b1;
        end else if (vmul_done) begin
            rd_reg <= {mul3_out, mul2_out, mul1_out, mul0_out};
            done   <= 1'b1;
        end else if (fmac_done) begin
            rd_reg <= {add3_out, add2_out, add1_out, add0_out};
            done   <= 1'b1;
        end else if (relu_done) begin
            rd_reg <= relu_result;
            done   <= 1'b1;
        end
    end
end

endmodule